/////////////////////***********************PACKAGE FOR PARAMETERS***********************/////////////////////
package mux_pkg;

  typedef struct {
    int WIDTH;
    int DEPTH;
    int SELECT_LINE_DEPTH;
  } mux_config_t;

endpackage
